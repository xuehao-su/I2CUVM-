
`define APB_DATA_WIDTH 32
`define APB_ADDR_WIDTH 32
